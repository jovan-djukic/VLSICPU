library verilog;
use verilog.vl_types.all;
entity SimpleInstructionTestBench is
    port(
        dummy           : in     vl_logic
    );
end SimpleInstructionTestBench;
