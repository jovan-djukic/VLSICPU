`ifndef SEVEN_SEGMENT_DISPLAY
`define SEVEN_SEGMENT_DISPLAY

`define ZERO		7'b1000000
`define ONE			7'b1111001
`define TWO			7'b0100100
`define THREE		7'b0110000
`define FOUR		7'b0011001
`define FIVE		7'b0010010
`define SIX			7'b0000010
`define SEVEN 		7'b1111000
`define EIGHT		7'b0000000
`define NINE		7'b0010000
`define TEN			7'b0001000
`define ELEVEN		7'b0000011
`define TWELVE		7'b1000110
`define THIRTEEN	7'b0100001
`define FOURTEEN	7'b0000100
`define FIFTEEN	7'b0001110

`define LOWER_ADDRESS	32'h2022
`define HIGHER_ADDRESS	32'h2023

`endif