`ifndef _TIMER_VH_
`define _TIMER_VH_

`timescale 1ps / 1ps

`endif