`ifndef _ALU_VH_
`define _ALU_VH_

`define ALU_ADD	0
`define ALU_SUB 1
`define ALU_MUL 2
`define ALU_DIV 3
`define ALU_SHR	4
`define ALU_SHL	5
`define ALU_AND	6
`define ALU_OR	7
`define ALU_NOT	8
`define ALU_A		9
`define	ALU_SWL	10
`define ALU_SWH	11
`define ALU_B 	12

`endif